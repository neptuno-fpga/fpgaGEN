package build_id is
constant BUILD_DATE : string := "201105";
constant BUILD_TIME : string := "123938";
end build_id;
