-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b80c3",
     9 => x"a8080b0b",
    10 => x"80c3ac08",
    11 => x"0b0b80c3",
    12 => x"b0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c3b00c0b",
    16 => x"0b80c3ac",
    17 => x"0c0b0b80",
    18 => x"c3a80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbbac",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c3a870",
    57 => x"80cde427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5190df",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c3",
    65 => x"b80c9f0b",
    66 => x"80c3bc0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c3bc08ff",
    70 => x"0580c3bc",
    71 => x"0c80c3bc",
    72 => x"088025e8",
    73 => x"3880c3b8",
    74 => x"08ff0580",
    75 => x"c3b80c80",
    76 => x"c3b80880",
    77 => x"25d03802",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"80c3b808",
    97 => x"25913882",
    98 => x"bc2d80c3",
    99 => x"b808ff05",
   100 => x"80c3b80c",
   101 => x"82fe0480",
   102 => x"c3b80880",
   103 => x"c3bc0853",
   104 => x"51728a2e",
   105 => x"098106be",
   106 => x"38715171",
   107 => x"9f24a438",
   108 => x"80c3b808",
   109 => x"a02911f8",
   110 => x"80115151",
   111 => x"a0713480",
   112 => x"c3bc0881",
   113 => x"0580c3bc",
   114 => x"0c80c3bc",
   115 => x"08519f71",
   116 => x"25de3880",
   117 => x"0b80c3bc",
   118 => x"0c80c3b8",
   119 => x"08810580",
   120 => x"c3b80c83",
   121 => x"fc0470a0",
   122 => x"2912f880",
   123 => x"11515172",
   124 => x"713480c3",
   125 => x"bc088105",
   126 => x"80c3bc0c",
   127 => x"80c3bc08",
   128 => x"a02e0981",
   129 => x"06913880",
   130 => x"0b80c3bc",
   131 => x"0c80c3b8",
   132 => x"08810580",
   133 => x"c3b80c02",
   134 => x"8c050d04",
   135 => x"02e8050d",
   136 => x"77795656",
   137 => x"880bfc16",
   138 => x"77712c8f",
   139 => x"06545254",
   140 => x"80537272",
   141 => x"25953871",
   142 => x"53fbe014",
   143 => x"51877134",
   144 => x"8114ff14",
   145 => x"545472f1",
   146 => x"387153f9",
   147 => x"1576712c",
   148 => x"87065351",
   149 => x"71802e8b",
   150 => x"38fbe014",
   151 => x"51717134",
   152 => x"81145472",
   153 => x"8e249538",
   154 => x"8f733153",
   155 => x"fbe01451",
   156 => x"a0713481",
   157 => x"14ff1454",
   158 => x"5472f138",
   159 => x"0298050d",
   160 => x"0402ec05",
   161 => x"0d800b80",
   162 => x"c3c00cf6",
   163 => x"8c08f690",
   164 => x"0871882c",
   165 => x"565481ff",
   166 => x"06527372",
   167 => x"25893871",
   168 => x"54820b80",
   169 => x"c3c00c72",
   170 => x"882c7381",
   171 => x"ff065455",
   172 => x"7473258d",
   173 => x"387280c3",
   174 => x"c0088407",
   175 => x"80c3c00c",
   176 => x"5573842b",
   177 => x"83f47125",
   178 => x"82713170",
   179 => x"0b0b0bbf",
   180 => x"940c8171",
   181 => x"2bf6880c",
   182 => x"fea413ff",
   183 => x"122c7888",
   184 => x"29ff9405",
   185 => x"70812c80",
   186 => x"c3c00852",
   187 => x"58525551",
   188 => x"52547680",
   189 => x"2e853870",
   190 => x"81075170",
   191 => x"f6940c71",
   192 => x"098105f6",
   193 => x"800c7209",
   194 => x"8105f684",
   195 => x"0c029405",
   196 => x"0d0402f4",
   197 => x"050d7453",
   198 => x"72708105",
   199 => x"5480f52d",
   200 => x"5271802e",
   201 => x"89387151",
   202 => x"82f82d86",
   203 => x"9804028c",
   204 => x"050d0402",
   205 => x"f4050d74",
   206 => x"70bfc206",
   207 => x"80cdc80c",
   208 => x"bfd07181",
   209 => x"06535353",
   210 => x"70881381",
   211 => x"b72d9812",
   212 => x"73822a70",
   213 => x"81065152",
   214 => x"52708813",
   215 => x"81b72d98",
   216 => x"1273832a",
   217 => x"70810651",
   218 => x"52527088",
   219 => x"1381b72d",
   220 => x"8c127384",
   221 => x"2a708106",
   222 => x"51525270",
   223 => x"881381b7",
   224 => x"2d72852a",
   225 => x"70810651",
   226 => x"53729413",
   227 => x"81b72d70",
   228 => x"80c3a80c",
   229 => x"028c050d",
   230 => x"0402f805",
   231 => x"0dbdac52",
   232 => x"80c3c451",
   233 => x"9fa62d80",
   234 => x"c3a80880",
   235 => x"2ea33880",
   236 => x"c6dc5280",
   237 => x"c3c451a1",
   238 => x"f32d80c6",
   239 => x"dc0880c3",
   240 => x"d00c80c6",
   241 => x"dc08fec0",
   242 => x"0c80c6dc",
   243 => x"085186b3",
   244 => x"2d028805",
   245 => x"0d0402f0",
   246 => x"050d8051",
   247 => x"94da2dbd",
   248 => x"ac5280c3",
   249 => x"c4519fa6",
   250 => x"2d80c3a8",
   251 => x"08802eaa",
   252 => x"3880c3d0",
   253 => x"0880c6dc",
   254 => x"0c80c6e0",
   255 => x"5480fd53",
   256 => x"80747084",
   257 => x"05560cff",
   258 => x"13537280",
   259 => x"25f23880",
   260 => x"c6dc5280",
   261 => x"c3c451a2",
   262 => x"9c2d0290",
   263 => x"050d0402",
   264 => x"d8050d80",
   265 => x"0bbfb40c",
   266 => x"80c3d008",
   267 => x"fec00c81",
   268 => x"0bfec40c",
   269 => x"840bfec4",
   270 => x"0c7b5280",
   271 => x"c3c4519f",
   272 => x"a62d80c3",
   273 => x"a8085380",
   274 => x"c3a80880",
   275 => x"2e818f38",
   276 => x"80c3c808",
   277 => x"57800bff",
   278 => x"18565874",
   279 => x"782e8b38",
   280 => x"81187581",
   281 => x"2a565874",
   282 => x"f738f718",
   283 => x"58815a80",
   284 => x"772580e3",
   285 => x"38775274",
   286 => x"51849c2d",
   287 => x"80c6dc52",
   288 => x"80c3c451",
   289 => x"a1f32d80",
   290 => x"c3a80880",
   291 => x"2ea83880",
   292 => x"c6dc5983",
   293 => x"fc567870",
   294 => x"84055a08",
   295 => x"7083ffff",
   296 => x"0671902a",
   297 => x"fec80cfe",
   298 => x"c80cfc17",
   299 => x"57537580",
   300 => x"25e43889",
   301 => x"be0480c3",
   302 => x"a8085a84",
   303 => x"805780c3",
   304 => x"c451a1c3",
   305 => x"2dfc8017",
   306 => x"81165657",
   307 => x"768024ff",
   308 => x"a4387980",
   309 => x"2e863882",
   310 => x"0bbfb40c",
   311 => x"79537280",
   312 => x"c3a80c02",
   313 => x"a8050d04",
   314 => x"02fc050d",
   315 => x"afc72dfe",
   316 => x"c4518171",
   317 => x"0c82710c",
   318 => x"0284050d",
   319 => x"0402f405",
   320 => x"0d747678",
   321 => x"53545280",
   322 => x"71259738",
   323 => x"72708105",
   324 => x"5480f52d",
   325 => x"72708105",
   326 => x"5481b72d",
   327 => x"ff115170",
   328 => x"eb388072",
   329 => x"81b72d02",
   330 => x"8c050d04",
   331 => x"02e8050d",
   332 => x"77568070",
   333 => x"56547376",
   334 => x"24b63880",
   335 => x"ccec0874",
   336 => x"2eae3873",
   337 => x"519ceb2d",
   338 => x"80c3a808",
   339 => x"80c3a808",
   340 => x"09810570",
   341 => x"80c3a808",
   342 => x"079f2a77",
   343 => x"05811757",
   344 => x"57535374",
   345 => x"76248938",
   346 => x"80ccec08",
   347 => x"7426d438",
   348 => x"7280c3a8",
   349 => x"0c029805",
   350 => x"0d0402f4",
   351 => x"050d80c2",
   352 => x"a4081551",
   353 => x"8aac2d80",
   354 => x"c3a80880",
   355 => x"2eac388b",
   356 => x"5380c3a8",
   357 => x"085280ca",
   358 => x"dc5189fd",
   359 => x"2d80cadc",
   360 => x"51889f2d",
   361 => x"80c3a808",
   362 => x"802e8f38",
   363 => x"bfb851b1",
   364 => x"ae2dafc7",
   365 => x"2d80518b",
   366 => x"c60480c2",
   367 => x"a851b1ae",
   368 => x"2dafb32d",
   369 => x"81518581",
   370 => x"2d028c05",
   371 => x"0d0402dc",
   372 => x"050d8070",
   373 => x"5a557480",
   374 => x"c2a40825",
   375 => x"b43880cc",
   376 => x"ec08752e",
   377 => x"ac387851",
   378 => x"9ceb2d80",
   379 => x"c3a80809",
   380 => x"81057080",
   381 => x"c3a80807",
   382 => x"9f2a7605",
   383 => x"811b5b56",
   384 => x"547480c2",
   385 => x"a4082589",
   386 => x"3880ccec",
   387 => x"087926d6",
   388 => x"38805578",
   389 => x"80ccec08",
   390 => x"2781db38",
   391 => x"78519ceb",
   392 => x"2d80c3a8",
   393 => x"08802e81",
   394 => x"ad3880c3",
   395 => x"a8088b05",
   396 => x"80f52d70",
   397 => x"842a7081",
   398 => x"06771078",
   399 => x"842b80ca",
   400 => x"dc0b80f5",
   401 => x"2d5c5c53",
   402 => x"51555673",
   403 => x"802e80cb",
   404 => x"38741682",
   405 => x"2b8e9a0b",
   406 => x"80c0f812",
   407 => x"0c547775",
   408 => x"311080c3",
   409 => x"d4115556",
   410 => x"90747081",
   411 => x"055681b7",
   412 => x"2da07481",
   413 => x"b72d7681",
   414 => x"ff068116",
   415 => x"58547380",
   416 => x"2e8a389c",
   417 => x"5380cadc",
   418 => x"528d9304",
   419 => x"8b5380c3",
   420 => x"a8085280",
   421 => x"c3d61651",
   422 => x"8dce0474",
   423 => x"16822b8a",
   424 => x"fa0b80c0",
   425 => x"f8120c54",
   426 => x"7681ff06",
   427 => x"81165854",
   428 => x"73802e8a",
   429 => x"389c5380",
   430 => x"cadc528d",
   431 => x"c5048b53",
   432 => x"80c3a808",
   433 => x"52777531",
   434 => x"1080c3d4",
   435 => x"05517655",
   436 => x"89fd2d8d",
   437 => x"eb047490",
   438 => x"29753170",
   439 => x"1080c3d4",
   440 => x"05515480",
   441 => x"c3a80874",
   442 => x"81b72d81",
   443 => x"1959748b",
   444 => x"24a3388c",
   445 => x"93047490",
   446 => x"29753170",
   447 => x"1080c3d4",
   448 => x"058c7731",
   449 => x"57515480",
   450 => x"7481b72d",
   451 => x"9e14ff16",
   452 => x"565474f3",
   453 => x"3802a405",
   454 => x"0d0402fc",
   455 => x"050d80c2",
   456 => x"a4081351",
   457 => x"8aac2d80",
   458 => x"c3a80880",
   459 => x"2e893880",
   460 => x"c3a80851",
   461 => x"94da2d80",
   462 => x"0b80c2a4",
   463 => x"0c8bce2d",
   464 => x"b08b2d02",
   465 => x"84050d04",
   466 => x"02fc050d",
   467 => x"725170fd",
   468 => x"2eb03870",
   469 => x"fd248a38",
   470 => x"70fc2e80",
   471 => x"cc388fb3",
   472 => x"0470fe2e",
   473 => x"b73870ff",
   474 => x"2e098106",
   475 => x"80c53880",
   476 => x"c2a40851",
   477 => x"70802ebb",
   478 => x"38ff1180",
   479 => x"c2a40c8f",
   480 => x"b30480c2",
   481 => x"a408f005",
   482 => x"7080c2a4",
   483 => x"0c517080",
   484 => x"25a13880",
   485 => x"0b80c2a4",
   486 => x"0c8fb304",
   487 => x"80c2a408",
   488 => x"810580c2",
   489 => x"a40c8fb3",
   490 => x"0480c2a4",
   491 => x"08900580",
   492 => x"c2a40c8b",
   493 => x"ce2db08b",
   494 => x"2d028405",
   495 => x"0d0402fc",
   496 => x"050d800b",
   497 => x"80c2a40c",
   498 => x"8bce2d80",
   499 => x"c0f051b1",
   500 => x"ae2d0284",
   501 => x"050d04bf",
   502 => x"fc0b80f5",
   503 => x"2d80c3a8",
   504 => x"0c0402fc",
   505 => x"050d7287",
   506 => x"065170bf",
   507 => x"fc0b81b7",
   508 => x"2d028405",
   509 => x"0d0402f8",
   510 => x"050d80cd",
   511 => x"c808bfc2",
   512 => x"06bfd80b",
   513 => x"80f52d52",
   514 => x"5270802e",
   515 => x"85387181",
   516 => x"0752bff0",
   517 => x"0b80f52d",
   518 => x"5170802e",
   519 => x"85387184",
   520 => x"075280c0",
   521 => x"880b80f5",
   522 => x"2d517080",
   523 => x"2e853871",
   524 => x"88075280",
   525 => x"c0940b80",
   526 => x"f52d5170",
   527 => x"802e8538",
   528 => x"71900752",
   529 => x"80c0a00b",
   530 => x"80f52d51",
   531 => x"70802e85",
   532 => x"3871a007",
   533 => x"527180c3",
   534 => x"a80c0288",
   535 => x"050d0402",
   536 => x"e0050d80",
   537 => x"0bbfb40c",
   538 => x"87558051",
   539 => x"86b32d74",
   540 => x"518fe22d",
   541 => x"810bfec4",
   542 => x"0c840bfe",
   543 => x"c40c830b",
   544 => x"fecc0cad",
   545 => x"802dafa7",
   546 => x"2dace32d",
   547 => x"ace32d81",
   548 => x"f92d8151",
   549 => x"85812dac",
   550 => x"e32dace3",
   551 => x"2d815185",
   552 => x"812dbdb8",
   553 => x"5186922d",
   554 => x"8453a6e2",
   555 => x"2d96802d",
   556 => x"80c3a808",
   557 => x"802e8638",
   558 => x"fe5391c5",
   559 => x"04ff1353",
   560 => x"728024e6",
   561 => x"3872802e",
   562 => x"82c03887",
   563 => x"992dbdd0",
   564 => x"51889f2d",
   565 => x"80c3a808",
   566 => x"802e9438",
   567 => x"bfb851b1",
   568 => x"ae2d8051",
   569 => x"85812d82",
   570 => x"0bbfb40c",
   571 => x"91fa0480",
   572 => x"c3a80851",
   573 => x"8fbe2daf",
   574 => x"b32dad99",
   575 => x"2db1c12d",
   576 => x"80c3a808",
   577 => x"80cdcc08",
   578 => x"882b80cd",
   579 => x"d00807fe",
   580 => x"d80c588f",
   581 => x"f62d80c3",
   582 => x"a80880c3",
   583 => x"d0082ea5",
   584 => x"3880c3a8",
   585 => x"0880c3d0",
   586 => x"0c80c3a8",
   587 => x"08fec00c",
   588 => x"84527751",
   589 => x"85812dac",
   590 => x"e32dace3",
   591 => x"2dff1252",
   592 => x"718025ee",
   593 => x"3880c054",
   594 => x"800bbf98",
   595 => x"57578653",
   596 => x"75708405",
   597 => x"570851ae",
   598 => x"e02d80c3",
   599 => x"a808812a",
   600 => x"70810651",
   601 => x"5271802e",
   602 => x"8d3880c3",
   603 => x"d0087432",
   604 => x"80c3d00c",
   605 => x"81577310",
   606 => x"ff145454",
   607 => x"728025d0",
   608 => x"38875376",
   609 => x"802e9038",
   610 => x"80c3d008",
   611 => x"fec00c80",
   612 => x"c3d00851",
   613 => x"86b32d85",
   614 => x"51aee02d",
   615 => x"80c3a808",
   616 => x"812a7081",
   617 => x"06515271",
   618 => x"802e9538",
   619 => x"ff157009",
   620 => x"709f2c72",
   621 => x"06705452",
   622 => x"53558fe2",
   623 => x"2db08b2d",
   624 => x"8651aee0",
   625 => x"2d80c3a8",
   626 => x"08812a70",
   627 => x"81065152",
   628 => x"71802e93",
   629 => x"38811555",
   630 => x"87752583",
   631 => x"38725574",
   632 => x"518fe22d",
   633 => x"b08b2d8f",
   634 => x"d72d80c3",
   635 => x"a808fed4",
   636 => x"0c77802e",
   637 => x"8c38bfb4",
   638 => x"088807fe",
   639 => x"c40c91fa",
   640 => x"04bfb408",
   641 => x"fec40c91",
   642 => x"fa04bddc",
   643 => x"5186922d",
   644 => x"800b80c3",
   645 => x"a80c02a0",
   646 => x"050d0402",
   647 => x"e8050d77",
   648 => x"797b5855",
   649 => x"55805372",
   650 => x"7625a338",
   651 => x"74708105",
   652 => x"5680f52d",
   653 => x"74708105",
   654 => x"5680f52d",
   655 => x"52527171",
   656 => x"2e863881",
   657 => x"5194d004",
   658 => x"81135394",
   659 => x"a7048051",
   660 => x"7080c3a8",
   661 => x"0c029805",
   662 => x"0d0402ec",
   663 => x"050d7655",
   664 => x"74802e80",
   665 => x"c2389a15",
   666 => x"80e02d51",
   667 => x"aba62d80",
   668 => x"c3a80880",
   669 => x"c3a80880",
   670 => x"cd8c0c80",
   671 => x"c3a80854",
   672 => x"5480cce8",
   673 => x"08802e9a",
   674 => x"38941580",
   675 => x"e02d51ab",
   676 => x"a62d80c3",
   677 => x"a808902b",
   678 => x"83fff00a",
   679 => x"06707507",
   680 => x"51537280",
   681 => x"cd8c0c80",
   682 => x"cd8c0853",
   683 => x"72802e9d",
   684 => x"3880cce0",
   685 => x"08fe1471",
   686 => x"2980ccf4",
   687 => x"080580cd",
   688 => x"900c7084",
   689 => x"2b80ccec",
   690 => x"0c5495fb",
   691 => x"0480ccf8",
   692 => x"0880cd8c",
   693 => x"0c80ccfc",
   694 => x"0880cd90",
   695 => x"0c80cce8",
   696 => x"08802e8b",
   697 => x"3880cce0",
   698 => x"08842b53",
   699 => x"95f60480",
   700 => x"cd800884",
   701 => x"2b537280",
   702 => x"ccec0c02",
   703 => x"94050d04",
   704 => x"02d8050d",
   705 => x"800b80cc",
   706 => x"e80c80c6",
   707 => x"dc528051",
   708 => x"a9d22d80",
   709 => x"c3a80854",
   710 => x"80c3a808",
   711 => x"8c38bdf0",
   712 => x"5186922d",
   713 => x"73559be8",
   714 => x"04805681",
   715 => x"0b80cd94",
   716 => x"0c8853bd",
   717 => x"fc5280c7",
   718 => x"9251949b",
   719 => x"2d80c3a8",
   720 => x"08762e09",
   721 => x"81068938",
   722 => x"80c3a808",
   723 => x"80cd940c",
   724 => x"8853be88",
   725 => x"5280c7ae",
   726 => x"51949b2d",
   727 => x"80c3a808",
   728 => x"893880c3",
   729 => x"a80880cd",
   730 => x"940c80cd",
   731 => x"9408802e",
   732 => x"81803880",
   733 => x"caa20b80",
   734 => x"f52d80ca",
   735 => x"a30b80f5",
   736 => x"2d71982b",
   737 => x"71902b07",
   738 => x"80caa40b",
   739 => x"80f52d70",
   740 => x"882b7207",
   741 => x"80caa50b",
   742 => x"80f52d71",
   743 => x"0780cada",
   744 => x"0b80f52d",
   745 => x"80cadb0b",
   746 => x"80f52d71",
   747 => x"882b0753",
   748 => x"5f54525a",
   749 => x"56575573",
   750 => x"81abaa2e",
   751 => x"0981068e",
   752 => x"387551aa",
   753 => x"f52d80c3",
   754 => x"a8085697",
   755 => x"db047382",
   756 => x"d4d52e87",
   757 => x"38be9451",
   758 => x"98a40480",
   759 => x"c6dc5275",
   760 => x"51a9d22d",
   761 => x"80c3a808",
   762 => x"5580c3a8",
   763 => x"08802e83",
   764 => x"f7388853",
   765 => x"be885280",
   766 => x"c7ae5194",
   767 => x"9b2d80c3",
   768 => x"a8088a38",
   769 => x"810b80cc",
   770 => x"e80c98aa",
   771 => x"048853bd",
   772 => x"fc5280c7",
   773 => x"9251949b",
   774 => x"2d80c3a8",
   775 => x"08802e8a",
   776 => x"38bea851",
   777 => x"86922d99",
   778 => x"890480ca",
   779 => x"da0b80f5",
   780 => x"2d547380",
   781 => x"d52e0981",
   782 => x"0680ce38",
   783 => x"80cadb0b",
   784 => x"80f52d54",
   785 => x"7381aa2e",
   786 => x"098106bd",
   787 => x"38800b80",
   788 => x"c6dc0b80",
   789 => x"f52d5654",
   790 => x"7481e92e",
   791 => x"83388154",
   792 => x"7481eb2e",
   793 => x"8c388055",
   794 => x"73752e09",
   795 => x"810682f8",
   796 => x"3880c6e7",
   797 => x"0b80f52d",
   798 => x"55748e38",
   799 => x"80c6e80b",
   800 => x"80f52d54",
   801 => x"73822e86",
   802 => x"3880559b",
   803 => x"e80480c6",
   804 => x"e90b80f5",
   805 => x"2d7080cc",
   806 => x"e00cff05",
   807 => x"80cce40c",
   808 => x"80c6ea0b",
   809 => x"80f52d80",
   810 => x"c6eb0b80",
   811 => x"f52d5876",
   812 => x"05778280",
   813 => x"29057080",
   814 => x"ccf00c80",
   815 => x"c6ec0b80",
   816 => x"f52d7080",
   817 => x"cd840c80",
   818 => x"cce80859",
   819 => x"57587680",
   820 => x"2e81b638",
   821 => x"8853be88",
   822 => x"5280c7ae",
   823 => x"51949b2d",
   824 => x"80c3a808",
   825 => x"82823880",
   826 => x"cce00870",
   827 => x"842b80cc",
   828 => x"ec0c7080",
   829 => x"cd800c80",
   830 => x"c7810b80",
   831 => x"f52d80c7",
   832 => x"800b80f5",
   833 => x"2d718280",
   834 => x"290580c7",
   835 => x"820b80f5",
   836 => x"2d708480",
   837 => x"80291280",
   838 => x"c7830b80",
   839 => x"f52d7081",
   840 => x"800a2912",
   841 => x"7080cd88",
   842 => x"0c80cd84",
   843 => x"08712980",
   844 => x"ccf00805",
   845 => x"7080ccf4",
   846 => x"0c80c789",
   847 => x"0b80f52d",
   848 => x"80c7880b",
   849 => x"80f52d71",
   850 => x"82802905",
   851 => x"80c78a0b",
   852 => x"80f52d70",
   853 => x"84808029",
   854 => x"1280c78b",
   855 => x"0b80f52d",
   856 => x"70982b81",
   857 => x"f00a0672",
   858 => x"057080cc",
   859 => x"f80cfe11",
   860 => x"7e297705",
   861 => x"80ccfc0c",
   862 => x"52595243",
   863 => x"545e5152",
   864 => x"59525d57",
   865 => x"59579be1",
   866 => x"0480c6ee",
   867 => x"0b80f52d",
   868 => x"80c6ed0b",
   869 => x"80f52d71",
   870 => x"82802905",
   871 => x"7080ccec",
   872 => x"0c70a029",
   873 => x"83ff0570",
   874 => x"892a7080",
   875 => x"cd800c80",
   876 => x"c6f30b80",
   877 => x"f52d80c6",
   878 => x"f20b80f5",
   879 => x"2d718280",
   880 => x"29057080",
   881 => x"cd880c7b",
   882 => x"71291e70",
   883 => x"80ccfc0c",
   884 => x"7d80ccf8",
   885 => x"0c730580",
   886 => x"ccf40c55",
   887 => x"5e515155",
   888 => x"55805194",
   889 => x"da2d8155",
   890 => x"7480c3a8",
   891 => x"0c02a805",
   892 => x"0d0402ec",
   893 => x"050d7670",
   894 => x"872c7180",
   895 => x"ff065556",
   896 => x"5480cce8",
   897 => x"088a3873",
   898 => x"882c7481",
   899 => x"ff065455",
   900 => x"80c6dc52",
   901 => x"80ccf008",
   902 => x"1551a9d2",
   903 => x"2d80c3a8",
   904 => x"085480c3",
   905 => x"a808802e",
   906 => x"b83880cc",
   907 => x"e808802e",
   908 => x"9a387284",
   909 => x"2980c6dc",
   910 => x"05700852",
   911 => x"53aaf52d",
   912 => x"80c3a808",
   913 => x"f00a0653",
   914 => x"9cdf0472",
   915 => x"1080c6dc",
   916 => x"057080e0",
   917 => x"2d5253ab",
   918 => x"a62d80c3",
   919 => x"a8085372",
   920 => x"547380c3",
   921 => x"a80c0294",
   922 => x"050d0402",
   923 => x"e0050d79",
   924 => x"70842c80",
   925 => x"cd900805",
   926 => x"718f0652",
   927 => x"5553728a",
   928 => x"3880c6dc",
   929 => x"527351a9",
   930 => x"d22d72a0",
   931 => x"2980c6dc",
   932 => x"05548074",
   933 => x"80f52d56",
   934 => x"5374732e",
   935 => x"83388153",
   936 => x"7481e52e",
   937 => x"81f43881",
   938 => x"70740654",
   939 => x"5872802e",
   940 => x"81e8388b",
   941 => x"1480f52d",
   942 => x"70832a79",
   943 => x"06585676",
   944 => x"9b3880c2",
   945 => x"d8085372",
   946 => x"89387280",
   947 => x"cadc0b81",
   948 => x"b72d7680",
   949 => x"c2d80c73",
   950 => x"539f9c04",
   951 => x"758f2e09",
   952 => x"810681b6",
   953 => x"38749f06",
   954 => x"8d2980ca",
   955 => x"cf115153",
   956 => x"811480f5",
   957 => x"2d737081",
   958 => x"055581b7",
   959 => x"2d831480",
   960 => x"f52d7370",
   961 => x"81055581",
   962 => x"b72d8514",
   963 => x"80f52d73",
   964 => x"70810555",
   965 => x"81b72d87",
   966 => x"1480f52d",
   967 => x"73708105",
   968 => x"5581b72d",
   969 => x"891480f5",
   970 => x"2d737081",
   971 => x"055581b7",
   972 => x"2d8e1480",
   973 => x"f52d7370",
   974 => x"81055581",
   975 => x"b72d9014",
   976 => x"80f52d73",
   977 => x"70810555",
   978 => x"81b72d92",
   979 => x"1480f52d",
   980 => x"73708105",
   981 => x"5581b72d",
   982 => x"941480f5",
   983 => x"2d737081",
   984 => x"055581b7",
   985 => x"2d961480",
   986 => x"f52d7370",
   987 => x"81055581",
   988 => x"b72d9814",
   989 => x"80f52d73",
   990 => x"70810555",
   991 => x"81b72d9c",
   992 => x"1480f52d",
   993 => x"73708105",
   994 => x"5581b72d",
   995 => x"9e1480f5",
   996 => x"2d7381b7",
   997 => x"2d7780c2",
   998 => x"d80c8053",
   999 => x"7280c3a8",
  1000 => x"0c02a005",
  1001 => x"0d0402cc",
  1002 => x"050d7e60",
  1003 => x"5e5a800b",
  1004 => x"80cd8c08",
  1005 => x"80cd9008",
  1006 => x"595c5680",
  1007 => x"5880ccec",
  1008 => x"08782e81",
  1009 => x"b838778f",
  1010 => x"06a01757",
  1011 => x"54739138",
  1012 => x"80c6dc52",
  1013 => x"76518117",
  1014 => x"57a9d22d",
  1015 => x"80c6dc56",
  1016 => x"807680f5",
  1017 => x"2d565474",
  1018 => x"742e8338",
  1019 => x"81547481",
  1020 => x"e52e80fd",
  1021 => x"38817075",
  1022 => x"06555c73",
  1023 => x"802e80f1",
  1024 => x"388b1680",
  1025 => x"f52d9806",
  1026 => x"597880e5",
  1027 => x"388b537c",
  1028 => x"52755194",
  1029 => x"9b2d80c3",
  1030 => x"a80880d5",
  1031 => x"389c1608",
  1032 => x"51aaf52d",
  1033 => x"80c3a808",
  1034 => x"841b0c9a",
  1035 => x"1680e02d",
  1036 => x"51aba62d",
  1037 => x"80c3a808",
  1038 => x"80c3a808",
  1039 => x"881c0c80",
  1040 => x"c3a80855",
  1041 => x"5580cce8",
  1042 => x"08802e99",
  1043 => x"38941680",
  1044 => x"e02d51ab",
  1045 => x"a62d80c3",
  1046 => x"a808902b",
  1047 => x"83fff00a",
  1048 => x"06701651",
  1049 => x"5473881b",
  1050 => x"0c787a0c",
  1051 => x"7b54a1b9",
  1052 => x"04811858",
  1053 => x"80ccec08",
  1054 => x"7826feca",
  1055 => x"3880cce8",
  1056 => x"08802eb3",
  1057 => x"387a519b",
  1058 => x"f22d80c3",
  1059 => x"a80880c3",
  1060 => x"a80880ff",
  1061 => x"fffff806",
  1062 => x"555b7380",
  1063 => x"fffffff8",
  1064 => x"2e953880",
  1065 => x"c3a808fe",
  1066 => x"0580cce0",
  1067 => x"082980cc",
  1068 => x"f4080557",
  1069 => x"9fbb0480",
  1070 => x"547380c3",
  1071 => x"a80c02b4",
  1072 => x"050d0402",
  1073 => x"f4050d74",
  1074 => x"70088105",
  1075 => x"710c7008",
  1076 => x"80cce408",
  1077 => x"06535371",
  1078 => x"8f388813",
  1079 => x"08519bf2",
  1080 => x"2d80c3a8",
  1081 => x"0888140c",
  1082 => x"810b80c3",
  1083 => x"a80c028c",
  1084 => x"050d0402",
  1085 => x"f0050d75",
  1086 => x"881108fe",
  1087 => x"0580cce0",
  1088 => x"082980cc",
  1089 => x"f4081172",
  1090 => x"0880cce4",
  1091 => x"08060579",
  1092 => x"55535454",
  1093 => x"a9d22d02",
  1094 => x"90050d04",
  1095 => x"02f0050d",
  1096 => x"75881108",
  1097 => x"fe0580cc",
  1098 => x"e0082980",
  1099 => x"ccf40811",
  1100 => x"720880cc",
  1101 => x"e4080605",
  1102 => x"79555354",
  1103 => x"54a8902d",
  1104 => x"0290050d",
  1105 => x"0402f405",
  1106 => x"0dd45281",
  1107 => x"ff720c71",
  1108 => x"085381ff",
  1109 => x"720c7288",
  1110 => x"2b83fe80",
  1111 => x"06720870",
  1112 => x"81ff0651",
  1113 => x"525381ff",
  1114 => x"720c7271",
  1115 => x"07882b72",
  1116 => x"087081ff",
  1117 => x"06515253",
  1118 => x"81ff720c",
  1119 => x"72710788",
  1120 => x"2b720870",
  1121 => x"81ff0672",
  1122 => x"0780c3a8",
  1123 => x"0c525302",
  1124 => x"8c050d04",
  1125 => x"02f4050d",
  1126 => x"74767181",
  1127 => x"ff06d40c",
  1128 => x"535380cd",
  1129 => x"98088538",
  1130 => x"71892b52",
  1131 => x"71982ad4",
  1132 => x"0c71902a",
  1133 => x"7081ff06",
  1134 => x"d40c5171",
  1135 => x"882a7081",
  1136 => x"ff06d40c",
  1137 => x"517181ff",
  1138 => x"06d40c72",
  1139 => x"902a7081",
  1140 => x"ff06d40c",
  1141 => x"51d40870",
  1142 => x"81ff0651",
  1143 => x"5182b8bf",
  1144 => x"527081ff",
  1145 => x"2e098106",
  1146 => x"943881ff",
  1147 => x"0bd40cd4",
  1148 => x"087081ff",
  1149 => x"06ff1454",
  1150 => x"515171e5",
  1151 => x"387080c3",
  1152 => x"a80c028c",
  1153 => x"050d0402",
  1154 => x"fc050d81",
  1155 => x"c75181ff",
  1156 => x"0bd40cff",
  1157 => x"11517080",
  1158 => x"25f43802",
  1159 => x"84050d04",
  1160 => x"02f0050d",
  1161 => x"a4872d8f",
  1162 => x"cf538052",
  1163 => x"87fc80f7",
  1164 => x"51a3942d",
  1165 => x"80c3a808",
  1166 => x"5480c3a8",
  1167 => x"08812e09",
  1168 => x"8106a438",
  1169 => x"81ff0bd4",
  1170 => x"0c820a52",
  1171 => x"849c80e9",
  1172 => x"51a3942d",
  1173 => x"80c3a808",
  1174 => x"8b3881ff",
  1175 => x"0bd40c73",
  1176 => x"53a4ee04",
  1177 => x"a4872dff",
  1178 => x"135372ff",
  1179 => x"bd387280",
  1180 => x"c3a80c02",
  1181 => x"90050d04",
  1182 => x"02f4050d",
  1183 => x"81ff0bd4",
  1184 => x"0c935380",
  1185 => x"5287fc80",
  1186 => x"c151a394",
  1187 => x"2d80c3a8",
  1188 => x"088b3881",
  1189 => x"ff0bd40c",
  1190 => x"8153a5a6",
  1191 => x"04a4872d",
  1192 => x"ff135372",
  1193 => x"de387280",
  1194 => x"c3a80c02",
  1195 => x"8c050d04",
  1196 => x"02f0050d",
  1197 => x"a4872d83",
  1198 => x"aa52849c",
  1199 => x"80c851a3",
  1200 => x"942d80c3",
  1201 => x"a808812e",
  1202 => x"09810693",
  1203 => x"38a2c52d",
  1204 => x"80c3a808",
  1205 => x"83ffff06",
  1206 => x"537283aa",
  1207 => x"2e9738a4",
  1208 => x"f82da5f0",
  1209 => x"048154a6",
  1210 => x"d804beb4",
  1211 => x"5186922d",
  1212 => x"8054a6d8",
  1213 => x"0481ff0b",
  1214 => x"d40cb153",
  1215 => x"a4a02d80",
  1216 => x"c3a80880",
  1217 => x"2e80c238",
  1218 => x"805287fc",
  1219 => x"80fa51a3",
  1220 => x"942d80c3",
  1221 => x"a808b238",
  1222 => x"81ff0bd4",
  1223 => x"0cd40853",
  1224 => x"81ff0bd4",
  1225 => x"0c81ff0b",
  1226 => x"d40c81ff",
  1227 => x"0bd40c81",
  1228 => x"ff0bd40c",
  1229 => x"72862a70",
  1230 => x"810680c3",
  1231 => x"a8085651",
  1232 => x"5372802e",
  1233 => x"9338a5e5",
  1234 => x"0472822e",
  1235 => x"ff9c38ff",
  1236 => x"135372ff",
  1237 => x"a7387254",
  1238 => x"7380c3a8",
  1239 => x"0c029005",
  1240 => x"0d0402f0",
  1241 => x"050d810b",
  1242 => x"80cd980c",
  1243 => x"8454d008",
  1244 => x"708f2a70",
  1245 => x"81065151",
  1246 => x"5372f338",
  1247 => x"72d00ca4",
  1248 => x"872dbec4",
  1249 => x"5186922d",
  1250 => x"d008708f",
  1251 => x"2a708106",
  1252 => x"51515372",
  1253 => x"f338810b",
  1254 => x"d00cb153",
  1255 => x"805284d4",
  1256 => x"80c051a3",
  1257 => x"942d80c3",
  1258 => x"a808812e",
  1259 => x"a1387282",
  1260 => x"2e098106",
  1261 => x"8c38bed0",
  1262 => x"5186922d",
  1263 => x"8053a886",
  1264 => x"04ff1353",
  1265 => x"72d638ff",
  1266 => x"145473ff",
  1267 => x"a138a5b0",
  1268 => x"2d80c3a8",
  1269 => x"0880cd98",
  1270 => x"0c80c3a8",
  1271 => x"088b3881",
  1272 => x"5287fc80",
  1273 => x"d051a394",
  1274 => x"2d81ff0b",
  1275 => x"d40cd008",
  1276 => x"708f2a70",
  1277 => x"81065151",
  1278 => x"5372f338",
  1279 => x"72d00c81",
  1280 => x"ff0bd40c",
  1281 => x"81537280",
  1282 => x"c3a80c02",
  1283 => x"90050d04",
  1284 => x"02e8050d",
  1285 => x"785681ff",
  1286 => x"0bd40cd0",
  1287 => x"08708f2a",
  1288 => x"70810651",
  1289 => x"515372f3",
  1290 => x"3882810b",
  1291 => x"d00c81ff",
  1292 => x"0bd40c77",
  1293 => x"5287fc80",
  1294 => x"d851a394",
  1295 => x"2d80c3a8",
  1296 => x"08802e8c",
  1297 => x"38bee851",
  1298 => x"86922d81",
  1299 => x"53a9c804",
  1300 => x"81ff0bd4",
  1301 => x"0c81fe0b",
  1302 => x"d40c80ff",
  1303 => x"55757084",
  1304 => x"05570870",
  1305 => x"982ad40c",
  1306 => x"70902c70",
  1307 => x"81ff06d4",
  1308 => x"0c547088",
  1309 => x"2c7081ff",
  1310 => x"06d40c54",
  1311 => x"7081ff06",
  1312 => x"d40c54ff",
  1313 => x"15557480",
  1314 => x"25d33881",
  1315 => x"ff0bd40c",
  1316 => x"81ff0bd4",
  1317 => x"0c81ff0b",
  1318 => x"d40c868d",
  1319 => x"a05481ff",
  1320 => x"0bd40cd4",
  1321 => x"0881ff06",
  1322 => x"55748738",
  1323 => x"ff145473",
  1324 => x"ed3881ff",
  1325 => x"0bd40cd0",
  1326 => x"08708f2a",
  1327 => x"70810651",
  1328 => x"515372f3",
  1329 => x"3872d00c",
  1330 => x"7280c3a8",
  1331 => x"0c029805",
  1332 => x"0d0402e8",
  1333 => x"050d7855",
  1334 => x"805681ff",
  1335 => x"0bd40cd0",
  1336 => x"08708f2a",
  1337 => x"70810651",
  1338 => x"515372f3",
  1339 => x"3882810b",
  1340 => x"d00c81ff",
  1341 => x"0bd40c77",
  1342 => x"5287fc80",
  1343 => x"d151a394",
  1344 => x"2d80dbc6",
  1345 => x"df5480c3",
  1346 => x"a808802e",
  1347 => x"8a38bef8",
  1348 => x"5186922d",
  1349 => x"aaeb0481",
  1350 => x"ff0bd40c",
  1351 => x"d4087081",
  1352 => x"ff065153",
  1353 => x"7281fe2e",
  1354 => x"0981069e",
  1355 => x"3880ff53",
  1356 => x"a2c52d80",
  1357 => x"c3a80875",
  1358 => x"70840557",
  1359 => x"0cff1353",
  1360 => x"728025ec",
  1361 => x"388156aa",
  1362 => x"d004ff14",
  1363 => x"5473c838",
  1364 => x"81ff0bd4",
  1365 => x"0c81ff0b",
  1366 => x"d40cd008",
  1367 => x"708f2a70",
  1368 => x"81065151",
  1369 => x"5372f338",
  1370 => x"72d00c75",
  1371 => x"80c3a80c",
  1372 => x"0298050d",
  1373 => x"0402f405",
  1374 => x"0d747088",
  1375 => x"2a83fe80",
  1376 => x"06707298",
  1377 => x"2a077288",
  1378 => x"2b87fc80",
  1379 => x"80067398",
  1380 => x"2b81f00a",
  1381 => x"06717307",
  1382 => x"0780c3a8",
  1383 => x"0c565153",
  1384 => x"51028c05",
  1385 => x"0d0402f8",
  1386 => x"050d028e",
  1387 => x"0580f52d",
  1388 => x"74882b07",
  1389 => x"7083ffff",
  1390 => x"0680c3a8",
  1391 => x"0c510288",
  1392 => x"050d0402",
  1393 => x"fc050d72",
  1394 => x"5180710c",
  1395 => x"800b8412",
  1396 => x"0c028405",
  1397 => x"0d0402f0",
  1398 => x"050d7570",
  1399 => x"08841208",
  1400 => x"535353ff",
  1401 => x"5471712e",
  1402 => x"a838afad",
  1403 => x"2d841308",
  1404 => x"70842914",
  1405 => x"88117008",
  1406 => x"7081ff06",
  1407 => x"84180881",
  1408 => x"11870684",
  1409 => x"1a0c5351",
  1410 => x"55515151",
  1411 => x"afa72d71",
  1412 => x"547380c3",
  1413 => x"a80c0290",
  1414 => x"050d0402",
  1415 => x"f8050daf",
  1416 => x"ad2de008",
  1417 => x"708b2a70",
  1418 => x"81065152",
  1419 => x"5270802e",
  1420 => x"a13880cd",
  1421 => x"9c087084",
  1422 => x"2980cda4",
  1423 => x"057381ff",
  1424 => x"06710c51",
  1425 => x"5180cd9c",
  1426 => x"08811187",
  1427 => x"0680cd9c",
  1428 => x"0c51800b",
  1429 => x"80cdc40c",
  1430 => x"af9f2daf",
  1431 => x"a72d0288",
  1432 => x"050d0402",
  1433 => x"fc050daf",
  1434 => x"ad2d810b",
  1435 => x"80cdc40c",
  1436 => x"afa72d80",
  1437 => x"cdc40851",
  1438 => x"70f93802",
  1439 => x"84050d04",
  1440 => x"02fc050d",
  1441 => x"80cd9c51",
  1442 => x"abc32dac",
  1443 => x"9b51af9b",
  1444 => x"2daec22d",
  1445 => x"0284050d",
  1446 => x"0402f405",
  1447 => x"0daea704",
  1448 => x"80c3a808",
  1449 => x"81f02e09",
  1450 => x"81068a38",
  1451 => x"810b80c3",
  1452 => x"9c0caea7",
  1453 => x"0480c3a8",
  1454 => x"0881e02e",
  1455 => x"0981068a",
  1456 => x"38810b80",
  1457 => x"c3a00cae",
  1458 => x"a70480c3",
  1459 => x"a8085280",
  1460 => x"c3a00880",
  1461 => x"2e893880",
  1462 => x"c3a80881",
  1463 => x"80055271",
  1464 => x"842c728f",
  1465 => x"06535380",
  1466 => x"c39c0880",
  1467 => x"2e9a3872",
  1468 => x"842980c2",
  1469 => x"dc057213",
  1470 => x"81712b70",
  1471 => x"09730806",
  1472 => x"730c5153",
  1473 => x"53ae9b04",
  1474 => x"72842980",
  1475 => x"c2dc0572",
  1476 => x"1383712b",
  1477 => x"72080772",
  1478 => x"0c535380",
  1479 => x"0b80c3a0",
  1480 => x"0c800b80",
  1481 => x"c39c0c80",
  1482 => x"cd9c51ab",
  1483 => x"d62d80c3",
  1484 => x"a808ff24",
  1485 => x"feea3880",
  1486 => x"0b80c3a8",
  1487 => x"0c028c05",
  1488 => x"0d0402f8",
  1489 => x"050d80c2",
  1490 => x"dc528f51",
  1491 => x"80727084",
  1492 => x"05540cff",
  1493 => x"11517080",
  1494 => x"25f23802",
  1495 => x"88050d04",
  1496 => x"02f0050d",
  1497 => x"7551afad",
  1498 => x"2d70822c",
  1499 => x"fc0680c2",
  1500 => x"dc117210",
  1501 => x"9e067108",
  1502 => x"70722a70",
  1503 => x"83068274",
  1504 => x"2b700974",
  1505 => x"06760c54",
  1506 => x"51565753",
  1507 => x"5153afa7",
  1508 => x"2d7180c3",
  1509 => x"a80c0290",
  1510 => x"050d0471",
  1511 => x"980c04ff",
  1512 => x"b00880c3",
  1513 => x"a80c0481",
  1514 => x"0bffb00c",
  1515 => x"04800bff",
  1516 => x"b00c0402",
  1517 => x"fc050d81",
  1518 => x"0b80c3a4",
  1519 => x"0c815185",
  1520 => x"812d0284",
  1521 => x"050d0402",
  1522 => x"fc050d80",
  1523 => x"0b80c3a4",
  1524 => x"0c805185",
  1525 => x"812d0284",
  1526 => x"050d0402",
  1527 => x"ec050d76",
  1528 => x"54805287",
  1529 => x"0b881580",
  1530 => x"f52d5653",
  1531 => x"74722483",
  1532 => x"38a05372",
  1533 => x"5182f82d",
  1534 => x"81128b15",
  1535 => x"80f52d54",
  1536 => x"52727225",
  1537 => x"de380294",
  1538 => x"050d0402",
  1539 => x"f0050d80",
  1540 => x"cdd40854",
  1541 => x"81f92d80",
  1542 => x"0b80cdd8",
  1543 => x"0c730880",
  1544 => x"2e818638",
  1545 => x"820b80c3",
  1546 => x"bc0c80cd",
  1547 => x"d8088f06",
  1548 => x"80c3b80c",
  1549 => x"73085271",
  1550 => x"832e9638",
  1551 => x"71832689",
  1552 => x"3871812e",
  1553 => x"af38b192",
  1554 => x"0471852e",
  1555 => x"9f38b192",
  1556 => x"04881480",
  1557 => x"f52d8415",
  1558 => x"08bf8853",
  1559 => x"54528692",
  1560 => x"2d718429",
  1561 => x"13700852",
  1562 => x"52b19604",
  1563 => x"7351afdb",
  1564 => x"2db19204",
  1565 => x"80cdc808",
  1566 => x"8815082c",
  1567 => x"70810651",
  1568 => x"5271802e",
  1569 => x"8738bf8c",
  1570 => x"51b18f04",
  1571 => x"bf905186",
  1572 => x"922d8414",
  1573 => x"08518692",
  1574 => x"2d80cdd8",
  1575 => x"08810580",
  1576 => x"cdd80c8c",
  1577 => x"1454b09d",
  1578 => x"04029005",
  1579 => x"0d047180",
  1580 => x"cdd40cb0",
  1581 => x"8b2d80cd",
  1582 => x"d808ff05",
  1583 => x"80cddc0c",
  1584 => x"0402e805",
  1585 => x"0d80cdd4",
  1586 => x"0880cde0",
  1587 => x"08575580",
  1588 => x"f851aee0",
  1589 => x"2d80c3a8",
  1590 => x"08812a70",
  1591 => x"81065152",
  1592 => x"719c3887",
  1593 => x"51aee02d",
  1594 => x"80c3a808",
  1595 => x"812a7081",
  1596 => x"06515271",
  1597 => x"802eb538",
  1598 => x"b1fe04ad",
  1599 => x"992d8751",
  1600 => x"aee02d80",
  1601 => x"c3a808f3",
  1602 => x"38b28f04",
  1603 => x"ad992d80",
  1604 => x"f851aee0",
  1605 => x"2d80c3a8",
  1606 => x"08f23880",
  1607 => x"c3a40881",
  1608 => x"327080c3",
  1609 => x"a40c7052",
  1610 => x"5285812d",
  1611 => x"800b80cd",
  1612 => x"cc0c800b",
  1613 => x"80cdd00c",
  1614 => x"80c3a408",
  1615 => x"838d3880",
  1616 => x"da51aee0",
  1617 => x"2d80c3a8",
  1618 => x"08802e8c",
  1619 => x"3880cdcc",
  1620 => x"08818007",
  1621 => x"80cdcc0c",
  1622 => x"80d951ae",
  1623 => x"e02d80c3",
  1624 => x"a808802e",
  1625 => x"8c3880cd",
  1626 => x"cc0880c0",
  1627 => x"0780cdcc",
  1628 => x"0c819451",
  1629 => x"aee02d80",
  1630 => x"c3a80880",
  1631 => x"2e8b3880",
  1632 => x"cdcc0890",
  1633 => x"0780cdcc",
  1634 => x"0c819151",
  1635 => x"aee02d80",
  1636 => x"c3a80880",
  1637 => x"2e8b3880",
  1638 => x"cdcc08a0",
  1639 => x"0780cdcc",
  1640 => x"0c81f551",
  1641 => x"aee02d80",
  1642 => x"c3a80880",
  1643 => x"2e8b3880",
  1644 => x"cdcc0881",
  1645 => x"0780cdcc",
  1646 => x"0c81f251",
  1647 => x"aee02d80",
  1648 => x"c3a80880",
  1649 => x"2e8b3880",
  1650 => x"cdcc0882",
  1651 => x"0780cdcc",
  1652 => x"0c81eb51",
  1653 => x"aee02d80",
  1654 => x"c3a80880",
  1655 => x"2e8b3880",
  1656 => x"cdcc0884",
  1657 => x"0780cdcc",
  1658 => x"0c81f451",
  1659 => x"aee02d80",
  1660 => x"c3a80880",
  1661 => x"2e8b3880",
  1662 => x"cdcc0888",
  1663 => x"0780cdcc",
  1664 => x"0c80d851",
  1665 => x"aee02d80",
  1666 => x"c3a80880",
  1667 => x"2e8c3880",
  1668 => x"cdd00881",
  1669 => x"800780cd",
  1670 => x"d00c9251",
  1671 => x"aee02d80",
  1672 => x"c3a80880",
  1673 => x"2e8c3880",
  1674 => x"cdd00880",
  1675 => x"c00780cd",
  1676 => x"d00c9451",
  1677 => x"aee02d80",
  1678 => x"c3a80880",
  1679 => x"2e8b3880",
  1680 => x"cdd00890",
  1681 => x"0780cdd0",
  1682 => x"0c9151ae",
  1683 => x"e02d80c3",
  1684 => x"a808802e",
  1685 => x"8b3880cd",
  1686 => x"d008a007",
  1687 => x"80cdd00c",
  1688 => x"9d51aee0",
  1689 => x"2d80c3a8",
  1690 => x"08802e8b",
  1691 => x"3880cdd0",
  1692 => x"08810780",
  1693 => x"cdd00c9b",
  1694 => x"51aee02d",
  1695 => x"80c3a808",
  1696 => x"802e8b38",
  1697 => x"80cdd008",
  1698 => x"820780cd",
  1699 => x"d00c9c51",
  1700 => x"aee02d80",
  1701 => x"c3a80880",
  1702 => x"2e8b3880",
  1703 => x"cdd00884",
  1704 => x"0780cdd0",
  1705 => x"0ca351ae",
  1706 => x"e02d80c3",
  1707 => x"a808802e",
  1708 => x"8b3880cd",
  1709 => x"d0088807",
  1710 => x"80cdd00c",
  1711 => x"81fd51ae",
  1712 => x"e02d81fa",
  1713 => x"51aee02d",
  1714 => x"bba00481",
  1715 => x"f551aee0",
  1716 => x"2d80c3a8",
  1717 => x"08812a70",
  1718 => x"81065152",
  1719 => x"71802eb3",
  1720 => x"3880cddc",
  1721 => x"08527180",
  1722 => x"2e8a38ff",
  1723 => x"1280cddc",
  1724 => x"0cb69304",
  1725 => x"80cdd808",
  1726 => x"1080cdd8",
  1727 => x"08057084",
  1728 => x"29165152",
  1729 => x"88120880",
  1730 => x"2e8938ff",
  1731 => x"51881208",
  1732 => x"52712d81",
  1733 => x"f251aee0",
  1734 => x"2d80c3a8",
  1735 => x"08812a70",
  1736 => x"81065152",
  1737 => x"71802eb4",
  1738 => x"3880cdd8",
  1739 => x"08ff1180",
  1740 => x"cddc0856",
  1741 => x"53537372",
  1742 => x"258a3881",
  1743 => x"1480cddc",
  1744 => x"0cb6dc04",
  1745 => x"72101370",
  1746 => x"84291651",
  1747 => x"52881208",
  1748 => x"802e8938",
  1749 => x"fe518812",
  1750 => x"0852712d",
  1751 => x"81fd51ae",
  1752 => x"e02d80c3",
  1753 => x"a808812a",
  1754 => x"70810651",
  1755 => x"5271802e",
  1756 => x"b13880cd",
  1757 => x"dc08802e",
  1758 => x"8a38800b",
  1759 => x"80cddc0c",
  1760 => x"b7a20480",
  1761 => x"cdd80810",
  1762 => x"80cdd808",
  1763 => x"05708429",
  1764 => x"16515288",
  1765 => x"1208802e",
  1766 => x"8938fd51",
  1767 => x"88120852",
  1768 => x"712d81fa",
  1769 => x"51aee02d",
  1770 => x"80c3a808",
  1771 => x"812a7081",
  1772 => x"06515271",
  1773 => x"802eb138",
  1774 => x"80cdd808",
  1775 => x"ff115452",
  1776 => x"80cddc08",
  1777 => x"73258938",
  1778 => x"7280cddc",
  1779 => x"0cb7e804",
  1780 => x"71101270",
  1781 => x"84291651",
  1782 => x"52881208",
  1783 => x"802e8938",
  1784 => x"fc518812",
  1785 => x"0852712d",
  1786 => x"80cddc08",
  1787 => x"70535473",
  1788 => x"802e8a38",
  1789 => x"8c15ff15",
  1790 => x"5555b7ef",
  1791 => x"04820b80",
  1792 => x"c3bc0c71",
  1793 => x"8f0680c3",
  1794 => x"b80c81eb",
  1795 => x"51aee02d",
  1796 => x"80c3a808",
  1797 => x"812a7081",
  1798 => x"06515271",
  1799 => x"802ead38",
  1800 => x"7408852e",
  1801 => x"098106a4",
  1802 => x"38881580",
  1803 => x"f52dff05",
  1804 => x"52718816",
  1805 => x"81b72d71",
  1806 => x"982b5271",
  1807 => x"80258838",
  1808 => x"800b8816",
  1809 => x"81b72d74",
  1810 => x"51afdb2d",
  1811 => x"81f451ae",
  1812 => x"e02d80c3",
  1813 => x"a808812a",
  1814 => x"70810651",
  1815 => x"5271802e",
  1816 => x"b3387408",
  1817 => x"852e0981",
  1818 => x"06aa3888",
  1819 => x"1580f52d",
  1820 => x"81055271",
  1821 => x"881681b7",
  1822 => x"2d7181ff",
  1823 => x"068b1680",
  1824 => x"f52d5452",
  1825 => x"72722787",
  1826 => x"38728816",
  1827 => x"81b72d74",
  1828 => x"51afdb2d",
  1829 => x"80da51ae",
  1830 => x"e02d80c3",
  1831 => x"a808812a",
  1832 => x"70810651",
  1833 => x"5271802e",
  1834 => x"81ad3880",
  1835 => x"cdd40880",
  1836 => x"cddc0855",
  1837 => x"5373802e",
  1838 => x"8a388c13",
  1839 => x"ff155553",
  1840 => x"b9b50472",
  1841 => x"08527182",
  1842 => x"2ea63871",
  1843 => x"82268938",
  1844 => x"71812eaa",
  1845 => x"38bad704",
  1846 => x"71832eb4",
  1847 => x"3871842e",
  1848 => x"09810680",
  1849 => x"f2388813",
  1850 => x"0851b1ae",
  1851 => x"2dbad704",
  1852 => x"80cddc08",
  1853 => x"51881308",
  1854 => x"52712dba",
  1855 => x"d704810b",
  1856 => x"8814082b",
  1857 => x"80cdc808",
  1858 => x"3280cdc8",
  1859 => x"0cbaab04",
  1860 => x"881380f5",
  1861 => x"2d81058b",
  1862 => x"1480f52d",
  1863 => x"53547174",
  1864 => x"24833880",
  1865 => x"54738814",
  1866 => x"81b72db0",
  1867 => x"8b2dbad7",
  1868 => x"04750880",
  1869 => x"2ea43875",
  1870 => x"0851aee0",
  1871 => x"2d80c3a8",
  1872 => x"08810652",
  1873 => x"71802e8c",
  1874 => x"3880cddc",
  1875 => x"08518416",
  1876 => x"0852712d",
  1877 => x"88165675",
  1878 => x"d8388054",
  1879 => x"800b80c3",
  1880 => x"bc0c738f",
  1881 => x"0680c3b8",
  1882 => x"0ca05273",
  1883 => x"80cddc08",
  1884 => x"2e098106",
  1885 => x"993880cd",
  1886 => x"d808ff05",
  1887 => x"74327009",
  1888 => x"81057072",
  1889 => x"079f2a91",
  1890 => x"71315151",
  1891 => x"53537151",
  1892 => x"82f82d81",
  1893 => x"14548e74",
  1894 => x"25c23880",
  1895 => x"c3a40852",
  1896 => x"7180c3a8",
  1897 => x"0c029805",
  1898 => x"0d040000",
  1899 => x"00ffffff",
  1900 => x"ff00ffff",
  1901 => x"ffff00ff",
  1902 => x"ffffff00",
  1903 => x"4f4b0000",
  1904 => x"52657365",
  1905 => x"74000000",
  1906 => x"53617665",
  1907 => x"20736574",
  1908 => x"74696e67",
  1909 => x"73000000",
  1910 => x"5363616e",
  1911 => x"6c696e65",
  1912 => x"73000000",
  1913 => x"41756469",
  1914 => x"6f20566f",
  1915 => x"6c756d65",
  1916 => x"00000000",
  1917 => x"4c6f6164",
  1918 => x"20524f4d",
  1919 => x"20100000",
  1920 => x"45786974",
  1921 => x"00000000",
  1922 => x"4d656761",
  1923 => x"64726976",
  1924 => x"65206d6f",
  1925 => x"64656c20",
  1926 => x"31000000",
  1927 => x"4d656761",
  1928 => x"64726976",
  1929 => x"65206d6f",
  1930 => x"64656c20",
  1931 => x"32000000",
  1932 => x"464d2064",
  1933 => x"69736162",
  1934 => x"6c650000",
  1935 => x"464d2065",
  1936 => x"6e61626c",
  1937 => x"65000000",
  1938 => x"50534720",
  1939 => x"64697361",
  1940 => x"626c6500",
  1941 => x"50534720",
  1942 => x"656e6162",
  1943 => x"6c650000",
  1944 => x"4a6f7973",
  1945 => x"7469636b",
  1946 => x"20737761",
  1947 => x"70000000",
  1948 => x"4a6f7973",
  1949 => x"7469636b",
  1950 => x"206e6f72",
  1951 => x"6d616c00",
  1952 => x"56474120",
  1953 => x"2d203331",
  1954 => x"4b487a00",
  1955 => x"5456202d",
  1956 => x"2031354b",
  1957 => x"487a0000",
  1958 => x"4261636b",
  1959 => x"00000000",
  1960 => x"4c6f6164",
  1961 => x"20457272",
  1962 => x"6f722100",
  1963 => x"46504741",
  1964 => x"47454e20",
  1965 => x"43464700",
  1966 => x"496e6974",
  1967 => x"69616c69",
  1968 => x"7a696e67",
  1969 => x"20534420",
  1970 => x"63617264",
  1971 => x"0a000000",
  1972 => x"424f4f54",
  1973 => x"20202020",
  1974 => x"47454e00",
  1975 => x"43617264",
  1976 => x"20696e69",
  1977 => x"74206661",
  1978 => x"696c6564",
  1979 => x"0a000000",
  1980 => x"4d425220",
  1981 => x"6661696c",
  1982 => x"0a000000",
  1983 => x"46415431",
  1984 => x"36202020",
  1985 => x"00000000",
  1986 => x"46415433",
  1987 => x"32202020",
  1988 => x"00000000",
  1989 => x"4e6f2070",
  1990 => x"61727469",
  1991 => x"74696f6e",
  1992 => x"20736967",
  1993 => x"0a000000",
  1994 => x"42616420",
  1995 => x"70617274",
  1996 => x"0a000000",
  1997 => x"53444843",
  1998 => x"20657272",
  1999 => x"6f72210a",
  2000 => x"00000000",
  2001 => x"53442069",
  2002 => x"6e69742e",
  2003 => x"2e2e0a00",
  2004 => x"53442063",
  2005 => x"61726420",
  2006 => x"72657365",
  2007 => x"74206661",
  2008 => x"696c6564",
  2009 => x"210a0000",
  2010 => x"57726974",
  2011 => x"65206661",
  2012 => x"696c6564",
  2013 => x"0a000000",
  2014 => x"52656164",
  2015 => x"20666169",
  2016 => x"6c65640a",
  2017 => x"00000000",
  2018 => x"16200000",
  2019 => x"14200000",
  2020 => x"15200000",
  2021 => x"00000002",
  2022 => x"00000016",
  2023 => x"0000001e",
  2024 => x"00000026",
  2025 => x"00000025",
  2026 => x"0000002e",
  2027 => x"00000036",
  2028 => x"0000003d",
  2029 => x"00000000",
  2030 => x"00000002",
  2031 => x"00001dc0",
  2032 => x"000004e8",
  2033 => x"00000002",
  2034 => x"00001dc8",
  2035 => x"000003d6",
  2036 => x"00000003",
  2037 => x"00002068",
  2038 => x"00000002",
  2039 => x"00000001",
  2040 => x"00001dd8",
  2041 => x"00000001",
  2042 => x"00000003",
  2043 => x"00002060",
  2044 => x"00000002",
  2045 => x"00000005",
  2046 => x"00001de4",
  2047 => x"00000007",
  2048 => x"00000003",
  2049 => x"00002058",
  2050 => x"00000002",
  2051 => x"00000003",
  2052 => x"00002050",
  2053 => x"00000002",
  2054 => x"00000003",
  2055 => x"00002048",
  2056 => x"00000002",
  2057 => x"00000002",
  2058 => x"00001df4",
  2059 => x"000007be",
  2060 => x"00000002",
  2061 => x"00001e00",
  2062 => x"000017c7",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00001e08",
  2067 => x"00001e1c",
  2068 => x"00001e30",
  2069 => x"00001e3c",
  2070 => x"00001e48",
  2071 => x"00001e54",
  2072 => x"00001e60",
  2073 => x"00001e70",
  2074 => x"00001e80",
  2075 => x"00001e8c",
  2076 => x"00000002",
  2077 => x"000021d4",
  2078 => x"0000057a",
  2079 => x"00000002",
  2080 => x"000021f2",
  2081 => x"0000057a",
  2082 => x"00000002",
  2083 => x"00002210",
  2084 => x"0000057a",
  2085 => x"00000002",
  2086 => x"0000222e",
  2087 => x"0000057a",
  2088 => x"00000002",
  2089 => x"0000224c",
  2090 => x"0000057a",
  2091 => x"00000002",
  2092 => x"0000226a",
  2093 => x"0000057a",
  2094 => x"00000002",
  2095 => x"00002288",
  2096 => x"0000057a",
  2097 => x"00000002",
  2098 => x"000022a6",
  2099 => x"0000057a",
  2100 => x"00000002",
  2101 => x"000022c4",
  2102 => x"0000057a",
  2103 => x"00000002",
  2104 => x"000022e2",
  2105 => x"0000057a",
  2106 => x"00000002",
  2107 => x"00002300",
  2108 => x"0000057a",
  2109 => x"00000002",
  2110 => x"0000231e",
  2111 => x"0000057a",
  2112 => x"00000002",
  2113 => x"0000233c",
  2114 => x"0000057a",
  2115 => x"00000004",
  2116 => x"00001e98",
  2117 => x"00001fb8",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000748",
  2121 => x"00000000",
  2122 => x"00000004",
  2123 => x"00001ea0",
  2124 => x"00001fb8",
  2125 => x"00000004",
  2126 => x"00001f40",
  2127 => x"00001fb8",
  2128 => x"00000004",
  2129 => x"00001dbc",
  2130 => x"00001fb8",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

