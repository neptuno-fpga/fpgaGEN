package build_id is
constant BUILD_DATE : string := "200424";
constant BUILD_TIME : string := "085604";
end build_id;
