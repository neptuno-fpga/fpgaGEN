package build_id is
constant BUILD_DATE : string := "201218";
constant BUILD_TIME : string := "214317";
end build_id;
