package build_id is
constant BUILD_DATE : string := "201004";
constant BUILD_TIME : string := "094433";
end build_id;
